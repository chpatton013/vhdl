package common is
  constant c_clock_rate: natural := 100000000; -- 100MHz
  constant c_clock_period: time := 1 sec / c_clock_rate;
end common;
